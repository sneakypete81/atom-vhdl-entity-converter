signal clk    : std_logic;
signal in     : std_logic_vector(WIDTH-1 downto 0);
signal output : std_logic_vector(WIDTH-1 downto 0);
