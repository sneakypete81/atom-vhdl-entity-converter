eNtiTy addWithCase Is
GeNeric (
  wiDTH  : Integer := 3;
  HEight : inTeger := 2
);
PorT (
  Clk    : In  STD_LOGIC;
  IN     : in  Std_Logic_Vector(width-1 DownTo 0);
  OutPut : oUt Std_Logic_Vector(width-1 DownTo 0)
);
EnD addWithCase;
