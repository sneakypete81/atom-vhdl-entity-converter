signal s_clk    : std_logic;
signal s_in     : std_logic_vector(WIDTH-1 downto 0);
signal s_output : std_logic_vector(WIDTH-1 downto 0);
