add_i : add
port map (
  clk    => clk,
  in     => in,
  output => output
);
